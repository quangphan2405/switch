package packet_pkg;
   
`include "packet_data.sv"   
`include "component_base.sv"
`include "sequencer.sv"
`include "monitor.sv"
`include "driver.sv"
`include "agent.sv"
`include "packet_vc.sv"

      
endpackage : packet_pkg
   
